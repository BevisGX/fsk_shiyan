library verilog;
use verilog.vl_types.all;
entity ENCODER is
    port(
        IN1             : in     vl_logic;
        IN2             : in     vl_logic;
        IN3             : in     vl_logic;
        IN4             : in     vl_logic;
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        \OUT\           : out    vl_logic
    );
end ENCODER;
